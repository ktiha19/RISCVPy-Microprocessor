module decoder();

endmodule